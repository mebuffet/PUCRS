
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41_USR5.90.69
#
# REF LIBS: lab3 
# TECH LIB NAME: cmos065
# TECH FILE NAME: techfile.cds
#******

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 1000  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;
LAYER PO
    TYPE MASTERSLICE ;
END PO

LAYER CO
    TYPE CUT ;
    SPACING 0.110 ;
    SPACING 0.140 ADJACENTCUTS 3 WITHIN 0.150 ;
END CO

LAYER M1
    TYPE ROUTING ;
    WIDTH 0.100 ;
    MINWIDTH 0.090 ;
    SPACING 0.090 ;
    OFFSET 0.000 ;
    PITCH 0.200 ;
    MINENCLOSEDAREA 0.200 ;
    DIRECTION VERTICAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 500.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 500.000 )  (  0.159 500.000 )  (  0.160 1000000.000 )  (  1.000 1000001.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO 5000.000 ;
    ANTENNACUMDIFFAREARATIO PWL  (  (  0.000 5000.000 )  (  0.159 5000.000 )  (  0.160 43072.960 )  (  1.000 43456.000 )  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END M1

LAYER VIA1
    TYPE CUT ;
    SPACING 0.100 ;
    SPACING 0.130 ADJACENTCUTS 3 WITHIN 0.140 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 20.000 )  (  0.159 20.000 )  (  0.160 933.600 )  (  1.000 1110.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFAREARATIO PWL  (  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END VIA1

LAYER M2
    TYPE ROUTING ;
    WIDTH 0.100 ;
    SPACING 0.100 ;
    OFFSET 0.000 ;
    PITCH 0.200 ;
    MINENCLOSEDAREA 0.200 ;
    DIRECTION HORIZONTAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 500.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 500.000 )  (  0.159 500.000 )  (  0.160 1000000.000 )  (  1.000 1000001.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO 5000.000 ;
    ANTENNACUMDIFFAREARATIO PWL  (  (  0.000 5000.000 )  (  0.159 5000.000 )  (  0.160 43072.960 )  (  1.000 43456.000 )  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END M2

LAYER VIA2
    TYPE CUT ;
    SPACING 0.100 ;
    SPACING 0.130 ADJACENTCUTS 3 WITHIN 0.140 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 20.000 )  (  0.159 20.000 )  (  0.160 933.600 )  (  1.000 1110.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFAREARATIO PWL  (  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END VIA2

LAYER M3
    TYPE ROUTING ;
    WIDTH 0.100 ;
    SPACING 0.100 ;
    OFFSET 0.000 ;
    PITCH 0.200 ;
    MINENCLOSEDAREA 0.200 ;
    DIRECTION VERTICAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 500.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 500.000 )  (  0.159 500.000 )  (  0.160 1000000.000 )  (  1.000 1000001.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO 5000.000 ;
    ANTENNACUMDIFFAREARATIO PWL  (  (  0.000 5000.000 )  (  0.159 5000.000 )  (  0.160 43072.960 )  (  1.000 43456.000 )  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END M3

LAYER VIA3
    TYPE CUT ;
    SPACING 0.100 ;
    SPACING 0.130 ADJACENTCUTS 3 WITHIN 0.140 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 20.000 )  (  0.159 20.000 )  (  0.160 933.600 )  (  1.000 1110.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFAREARATIO PWL  (  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END VIA3

LAYER M4
    TYPE ROUTING ;
    WIDTH 0.100 ;
    SPACING 0.100 ;
    OFFSET 0.000 ;
    PITCH 0.200 ;
    MINENCLOSEDAREA 0.200 ;
    DIRECTION HORIZONTAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 500.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 500.000 )  (  0.159 500.000 )  (  0.160 1000000.000 )  (  1.000 1000001.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO 5000.000 ;
    ANTENNACUMDIFFAREARATIO PWL  (  (  0.000 5000.000 )  (  0.159 5000.000 )  (  0.160 43072.960 )  (  1.000 43456.000 )  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END M4

LAYER VIA4
    TYPE CUT ;
    SPACING 0.100 ;
    SPACING 0.130 ADJACENTCUTS 3 WITHIN 0.140 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 20.000 )  (  0.159 20.000 )  (  0.160 933.600 )  (  1.000 1110.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFAREARATIO PWL  (  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END VIA4

LAYER M5
    TYPE ROUTING ;
    WIDTH 0.100 ;
    SPACING 0.100 ;
    OFFSET 0.000 ;
    PITCH 0.200 ;
    MINENCLOSEDAREA 0.200 ;
    DIRECTION VERTICAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 500.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 500.000 )  (  0.159 500.000 )  (  0.160 1000000.000 )  (  1.000 1000001.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO 5000.000 ;
    ANTENNACUMDIFFAREARATIO PWL  (  (  0.000 5000.000 )  (  0.159 5000.000 )  (  0.160 43072.960 )  (  1.000 43456.000 )  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END M5

LAYER VIA5
    TYPE CUT ;
    SPACING 0.540 ;
    SPACING 0.540 ADJACENTCUTS 3 WITHIN 0.560 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 20.000 )  (  0.159 20.000 )  (  0.160 933.600 )  (  1.000 1110.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFAREARATIO PWL  (  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END VIA5

LAYER M6
    TYPE ROUTING ;
    WIDTH 0.400 ;
    SPACING 0.400 ;
    OFFSET 0.000 ;
    PITCH 0.800 ;
    MINENCLOSEDAREA 0.565 ;
    DIRECTION HORIZONTAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 500.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 500.000 )  (  0.159 500.000 )  (  0.160 1000000.000 )  (  1.000 1000001.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO 5000.000 ;
    ANTENNACUMDIFFAREARATIO PWL  (  (  0.000 5000.000 )  (  0.159 5000.000 )  (  0.160 43072.960 )  (  1.000 43456.000 )  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END M6

LAYER VIA6
    TYPE CUT ;
    SPACING 0.540 ;
    SPACING 0.540 ADJACENTCUTS 3 WITHIN 0.560 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 20.000 )  (  0.159 20.000 )  (  0.160 933.600 )  (  1.000 1110.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFAREARATIO PWL  (  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END VIA6

LAYER M7
    TYPE ROUTING ;
    WIDTH 0.400 ;
    SPACING 0.400 ;
    OFFSET 0.000 ;
    PITCH 0.800 ;
    MINENCLOSEDAREA 0.565 ;
    DIRECTION VERTICAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 500.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 500.000 )  (  0.159 500.000 )  (  0.160 1000000.000 )  (  1.000 1000001.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO 5000.000 ;
    ANTENNACUMDIFFAREARATIO PWL  (  (  0.000 5000.000 )  (  0.159 5000.000 )  (  0.160 43072.960 )  (  1.000 43456.000 )  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END M7

LAYER CB
    TYPE CUT ;
    SPACING 2.000 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 20.000 )  (  0.159 20.000 )  (  0.160 933.600 )  (  1.000 1110.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFAREARATIO PWL  (  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END CB

LAYER AP
    TYPE ROUTING ;
    WIDTH 3.000 ;
    SPACING 2.000 ;
    OFFSET 0.000 ;
    PITCH 5.000 ;
    DIRECTION HORIZONTAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 500.000 ;
    ANTENNASIDEAREARATIO PWL  (  )  ;
    ANTENNADIFFAREARATIO PWL  (  (  0.000 500.000 )  (  0.159 500.000 )  (  0.160 1000000.000 )  (  1.000 1000001.000 )  )  ;
    ANTENNADIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMAREARATIO 5000.000 ;
    ANTENNACUMDIFFAREARATIO PWL  (  (  0.000 5000.000 )  (  0.159 5000.000 )  (  0.160 43072.960 )  (  1.000 43456.000 )  )  ;
    ANTENNACUMSIDEAREARATIO PWL  (  )  ;
    ANTENNACUMDIFFSIDEAREARATIO PWL  (  )  ;
    ANTENNAAREAFACTOR  ;
    ANTENNASIDEAREAFACTOR  ;
END AP

LAYER overlap
    TYPE OVERLAP ;
END overlap

VIA PTAP_
    LAYER M1 ;
        RECT -0.045 -0.085 0.045 0.085 ;
    LAYER CO ;
        RECT -0.045 -0.045 0.045 0.045 ;
    LAYER PP ;
        RECT -0.095 -0.095 0.095 0.095 ;
END PTAP_

VIA NTAP_
    LAYER M1 ;
        RECT -0.045 -0.085 0.045 0.085 ;
    LAYER CO ;
        RECT -0.045 -0.045 0.045 0.045 ;
    LAYER NP ;
        RECT -0.095 -0.095 0.095 0.095 ;
END NTAP_

VIA M1__POD
    LAYER M1 ;
        RECT -0.045 -0.085 0.045 0.085 ;
    LAYER CO ;
        RECT -0.045 -0.045 0.045 0.045 ;
    LAYER OD ;
        RECT -0.075 -0.075 0.075 0.075 ;
END M1__POD

VIA M1__NOD
    LAYER M1 ;
        RECT -0.045 -0.085 0.045 0.085 ;
    LAYER CO ;
        RECT -0.045 -0.045 0.045 0.045 ;
    LAYER OD ;
        RECT -0.075 -0.075 0.075 0.075 ;
END M1__NOD

VIA M1__NW
    LAYER M1 ;
        RECT -0.045 -0.085 0.045 0.085 ;
    LAYER CO ;
        RECT -0.045 -0.045 0.045 0.045 ;
    LAYER NW ;
        RECT -0.235 -0.235 0.235 0.235 ;
END M1__NW

VIA M1__OD
    LAYER M1 ;
        RECT -0.045 -0.085 0.045 0.085 ;
    LAYER CO ;
        RECT -0.045 -0.045 0.045 0.045 ;
    LAYER OD ;
        RECT -0.075 -0.075 0.075 0.075 ;
END M1__OD

VIA M2X_PO
    LAYER M2 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER PO ;
        RECT -0.055 -0.085 0.055 0.085 ;
END M2X_PO

VIA M3X_PO
    LAYER M3 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER PO ;
        RECT -0.055 -0.085 0.055 0.085 ;
END M3X_PO

VIA M3X_M1
    LAYER M3 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M1 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M3X_M1

VIA M4X_PO
    LAYER M4 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER PO ;
        RECT -0.055 -0.085 0.055 0.085 ;
END M4X_PO

VIA M4X_M1
    LAYER M4 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M1 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M4X_M1

VIA M4X_M2X
    LAYER M4 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M4X_M2X

VIA M5X_PO
    LAYER M5 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER PO ;
        RECT -0.055 -0.085 0.055 0.085 ;
END M5X_PO

VIA M5X_M1
    LAYER M5 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M1 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M5X_M1

VIA M5X_M2X
    LAYER M5 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M5X_M2X

VIA M5X_M3X
    LAYER M5 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M3 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M5X_M3X

VIA M6Z_PO
    LAYER PO ;
        RECT -0.055 -0.085 0.055 0.085 ;
END M6Z_PO

VIA M6Z_M1
    LAYER M1 ;
        RECT -0.150 -0.190 0.150 0.190 ;
END M6Z_M1

VIA M6Z_M2X
    LAYER M2 ;
        RECT -0.150 -0.190 0.150 0.190 ;
END M6Z_M2X

VIA M6Z_M3X
    LAYER M3 ;
        RECT -0.150 -0.190 0.150 0.190 ;
END M6Z_M3X

VIA M6Z_M4X
    LAYER M4 ;
        RECT -0.150 -0.190 0.150 0.190 ;
END M6Z_M4X

VIA M7Z_PO
    LAYER PO ;
        RECT -0.055 -0.085 0.055 0.085 ;
END M7Z_PO

VIA M7Z_M1
    LAYER M1 ;
        RECT -0.150 -0.190 0.150 0.190 ;
END M7Z_M1

VIA M7Z_M2X
    LAYER M2 ;
        RECT -0.150 -0.190 0.150 0.190 ;
END M7Z_M2X

VIA M7Z_M3X
    LAYER M3 ;
        RECT -0.150 -0.190 0.150 0.190 ;
END M7Z_M3X

VIA M7Z_M4X
    LAYER M4 ;
        RECT -0.150 -0.190 0.150 0.190 ;
END M7Z_M4X

VIA M7Z_M5X
    LAYER M5 ;
        RECT -0.200 -0.260 0.200 0.260 ;
END M7Z_M5X

VIA M1__PO
    LAYER PO ;
        RECT -0.055 -0.085 0.055 0.085 ;
    LAYER CO ;
        RECT -0.045 -0.045 0.045 0.045 ;
    LAYER M1 ;
        RECT -0.085 -0.045 0.085 0.045 ;
END M1__PO

VIA M2X_M1 DEFAULT
    LAYER M1 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M2X_M1

VIA M2X_M1_H DEFAULT
    LAYER M1 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M2 ;
        RECT -0.090 -0.050 0.090 0.050 ;
END M2X_M1_H

VIA M2X_M1_V
    LAYER M1 ;
        RECT -0.090 -0.050 0.090 0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M2X_M1_V

VIA M3X_M2X DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M3 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M3X_M2X

VIA M3X_M2X_H DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050 0.090 0.050 ;
END M3X_M2X_H

VIA M3X_M2X_V
    LAYER M2 ;
        RECT -0.090 -0.050 0.090 0.050 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M3 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M3X_M2X_V

VIA M4X_M3X DEFAULT
    LAYER M3 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M4X_M3X

VIA M4X_M3X_H DEFAULT
    LAYER M3 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M4 ;
        RECT -0.090 -0.050 0.090 0.050 ;
END M4X_M3X_H

VIA M4X_M3X_V
    LAYER M3 ;
        RECT -0.090 -0.050 0.090 0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M4X_M3X_V

VIA M5X_M4X DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M5 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M5X_M4X

VIA M5X_M4X_H DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.090 0.050 0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050 0.090 0.050 ;
END M5X_M4X_H

VIA M5X_M4X_V
    LAYER M4 ;
        RECT -0.090 -0.050 0.090 0.050 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050 0.050 0.050 ;
    LAYER M5 ;
        RECT -0.050 -0.090 0.050 0.090 ;
END M5X_M4X_V

VIA M6Z__M5X DEFAULT
    LAYER M5 ;
        RECT -0.200 -0.260 0.200 0.260 ;
END M6Z__M5X

VIA M6Z__M5X_H DEFAULT
    LAYER M5 ;
        RECT -0.200 -0.260 0.200 0.260 ;
END M6Z__M5X_H

VIA M6Z_M5X_V
    LAYER M5 ;
        RECT -0.260 -0.200 0.260 0.200 ;
END M6Z_M5X_V

VIA M7Z__M6Z DEFAULT
END M7Z__M6Z

VIA M7Z__M6Z_H DEFAULT
END M7Z__M6Z_H

VIA M7Z_M6Z_V
END M7Z_M6Z_V

VIA AP__M7Z DEFAULT
    LAYER CB ;
        RECT -1.500 -1.500 1.500 1.500 ;
    LAYER AP ;
        RECT -2.200 -2.200 2.200 2.200 ;
END AP__M7Z

VIA M6Z__BOTMIM
    LAYER BOTMIM ;
        RECT -0.780 -0.780 0.780 0.780 ;
END M6Z__BOTMIM

VIA M6Z__MKTOPMIM
    LAYER MKTOPMIM ;
        RECT -0.780 -0.780 0.780 0.780 ;
END M6Z__MKTOPMIM

SITE CoreSite
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.200 BY 2.600 ;
END CoreSite

MACRO Complex_f2
    CLASS CORE ;
    FOREIGN Complex_f2 0 -2.8 ;
    ORIGIN 0.000 2.800 ;
    SIZE 2.200 BY 2.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.605 -1.215 0.755 -0.815 ;
        RECT  0.605 -1.395 0.695 -0.815 ;
        RECT  0.230 -1.395 0.695 -1.305 ;
        RECT  0.230 -2.185 0.380 -1.805 ;
        RECT  0.230 -2.185 0.320 -1.305 ;
        END
    END S
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 -1.700 2.000 -1.550 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -1.700 1.580 -1.550 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 -1.700 1.160 -1.550 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 -1.700 0.740 -1.550 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.560 2.200 0.000 ;
        RECT  1.820 -1.215 1.970 -0.815 ;
        RECT  1.850 -1.215 1.940 0.000 ;
        RECT  0.230 -1.215 0.380 -0.815 ;
        RECT  0.260 -1.215 0.350 0.000 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -3.000 2.200 -2.440 ;
        RECT  1.820 -2.185 1.970 -1.985 ;
        RECT  1.850 -3.000 1.940 -1.985 ;
        RECT  1.025 -2.185 1.175 -1.985 ;
        RECT  1.055 -3.000 1.145 -1.985 ;
        END
    END gnd!
    OBS
        LAYER M1 ;
        RECT  0.605 -2.185 0.755 -1.985 ;
        RECT  1.445 -2.185 1.595 -1.985 ;
        RECT  0.665 -2.185 0.755 -1.805 ;
        RECT  1.445 -2.185 1.535 -1.805 ;
        RECT  0.665 -1.895 1.535 -1.805 ;
    END
END Complex_f2

END LIBRARY
