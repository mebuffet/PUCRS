
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41_USR5.90.69
#
# REF LIBS: lab3 
# TECH LIB NAME: cmos065
# TECH FILE NAME: techfile.cds
#******

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 1000  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;
SITE CORE
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.200 BY 2.600 ;
END CORE

MACRO Complex_f2
    CLASS CORE ;
    FOREIGN Complex_f2 0 -2.8 ;
    ORIGIN 0.000 2.800 ;
    SIZE 2.200 BY 2.600 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.025 -1.215 1.175 -0.815 ;
        RECT  1.025 -1.395 1.115 -0.815 ;
        RECT  0.290 -1.395 1.115 -1.305 ;
        RECT  0.635 -1.895 0.725 -1.305 ;
        RECT  0.230 -1.895 0.725 -1.805 ;
        RECT  0.230 -1.215 0.380 -0.815 ;
        RECT  0.290 -1.395 0.380 -0.815 ;
        RECT  0.230 -2.185 0.380 -1.805 ;
        END
    END S
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 -1.700 2.000 -1.550 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -1.700 1.580 -1.550 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 -1.700 1.160 -1.550 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 -1.700 0.500 -1.550 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.560 2.200 0.000 ;
        RECT  1.880 -1.215 1.970 0.000 ;
        RECT  1.820 -1.215 1.970 -0.815 ;
        RECT  0.605 -1.215 0.755 -0.815 ;
        RECT  0.635 -1.215 0.725 0.000 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -3.000 2.200 -2.440 ;
        RECT  1.445 -2.185 1.595 -1.985 ;
        RECT  1.475 -3.000 1.565 -1.985 ;
        END
    END gnd!
    OBS
        LAYER M1 ;
        RECT  1.025 -2.185 1.175 -1.985 ;
        RECT  1.820 -2.185 1.970 -1.985 ;
        RECT  1.085 -2.185 1.175 -1.805 ;
        RECT  1.820 -2.185 1.910 -1.805 ;
        RECT  1.085 -1.895 1.910 -1.805 ;
    END
END Complex_f2

END LIBRARY
